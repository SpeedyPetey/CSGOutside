// ============================================================================
// Copyright (c) 2013 by Terasic Technologies Inc.
// ============================================================================
//
// Permission:
//
//   Terasic grants permission to use and modify this code for use
//   in synthesis for all Terasic Development Boards and Altera Development 
//   Kits made by Terasic.  Other use of this code, including the selling 
//   ,duplication, or modification of any portion is strictly prohibited.
//
// Disclaimer:
//
//   This VHDL/Verilog or C/C++ source code is intended as a design reference
//   which illustrates how these types of functions can be implemented.
//   It is the user's responsibility to verify their design for
//   consistency and functionality through the use of formal
//   verification methods.  Terasic provides no warranty regarding the use 
//   or functionality of this code.
//
// ============================================================================
//           
//  Terasic Technologies Inc
//  9F., No.176, Sec.2, Gongdao 5th Rd, East Dist, Hsinchu City, 30070. Taiwan
//  
//  
//                     web: http://www.terasic.com/  
//                     email: support@terasic.com
//
// ============================================================================
//Date:  Mon Jun 17 20:35:29 2013
// ============================================================================

//`define ENABLE_HPS

module DE1_SoC_Audio(

      ///////// ADC /////////
      output             ADC_CONVST,
      output             ADC_DIN,
      input              ADC_DOUT,
      output             ADC_SCLK,

      ///////// AUD /////////
      input              AUD_ADCDAT,
      inout              AUD_ADCLRCK,
      inout              AUD_BCLK,
      output             AUD_DACDAT,
      inout              AUD_DACLRCK,
      output             AUD_XCK,

      ///////// CLOCK2 /////////
      input              CLOCK2_50,

      ///////// CLOCK3 /////////
      input              CLOCK3_50,

      ///////// CLOCK4 /////////
      input              CLOCK4_50,

      ///////// CLOCK /////////
      input              CLOCK_50,

      ///////// DRAM /////////
      output      [12:0] DRAM_ADDR,
      output      [1:0]  DRAM_BA,
      output             DRAM_CAS_N,
      output             DRAM_CKE,
      output             DRAM_CLK,
      output             DRAM_CS_N,
      inout       [15:0] DRAM_DQ,
      output             DRAM_LDQM,
      output             DRAM_RAS_N,
      output             DRAM_UDQM,
      output             DRAM_WE_N,

      ///////// FAN /////////
      output             FAN_CTRL,

      ///////// FPGA /////////
      output             FPGA_I2C_SCLK,
      inout              FPGA_I2C_SDAT,

      ///////// GPIO /////////
      inout     [35:0]         GPIO_0,
      inout     [35:0]         GPIO_1,
 


`ifdef ENABLE_HPS
      ///////// HPS /////////
      inout              HPS_CONV_USB_N,
      output      [14:0] HPS_DDR3_ADDR,
      output      [2:0]  HPS_DDR3_BA,
      output             HPS_DDR3_CAS_N,
      output             HPS_DDR3_CKE,
      output             HPS_DDR3_CK_N,
      output             HPS_DDR3_CK_P,
      output             HPS_DDR3_CS_N,
      output      [3:0]  HPS_DDR3_DM,
      inout       [31:0] HPS_DDR3_DQ,
      inout       [3:0]  HPS_DDR3_DQS_N,
      inout       [3:0]  HPS_DDR3_DQS_P,
      output             HPS_DDR3_ODT,
      output             HPS_DDR3_RAS_N,
      output             HPS_DDR3_RESET_N,
      input              HPS_DDR3_RZQ,
      output             HPS_DDR3_WE_N,
      output             HPS_ENET_GTX_CLK,
      inout              HPS_ENET_INT_N,
      output             HPS_ENET_MDC,
      inout              HPS_ENET_MDIO,
      input              HPS_ENET_RX_CLK,
      input       [3:0]  HPS_ENET_RX_DATA,
      input              HPS_ENET_RX_DV,
      output      [3:0]  HPS_ENET_TX_DATA,
      output             HPS_ENET_TX_EN,
      inout       [3:0]  HPS_FLASH_DATA,
      output             HPS_FLASH_DCLK,
      output             HPS_FLASH_NCSO,
      inout              HPS_GSENSOR_INT,
      inout              HPS_I2C1_SCLK,
      inout              HPS_I2C1_SDAT,
      inout              HPS_I2C2_SCLK,
      inout              HPS_I2C2_SDAT,
      inout              HPS_I2C_CONTROL,
      inout              HPS_KEY,
      inout              HPS_LED,
      inout              HPS_LTC_GPIO,
      output             HPS_SD_CLK,
      inout              HPS_SD_CMD,
      inout       [3:0]  HPS_SD_DATA,
      output             HPS_SPIM_CLK,
      input              HPS_SPIM_MISO,
      output             HPS_SPIM_MOSI,
      inout              HPS_SPIM_SS,
      input              HPS_UART_RX,
      output             HPS_UART_TX,
      input              HPS_USB_CLKOUT,
      inout       [7:0]  HPS_USB_DATA,
      input              HPS_USB_DIR,
      input              HPS_USB_NXT,
      output             HPS_USB_STP,
`endif /*ENABLE_HPS*/

      ///////// IRDA /////////
      input              IRDA_RXD,
      output             IRDA_TXD,

		input [3:0] KEY,
		output [6:0] HEX0, output [6:0] HEX1, output [6:0] HEX2,
      //output [6:0] HEX3, output [6:0] HEX4, output [6:0] HEX5,
		output [9:0] LEDR,

      ///////// PS2 /////////
      inout              PS2_CLK,
      inout              PS2_CLK2,
      inout              PS2_DAT,
      inout              PS2_DAT2,

      ///////// TD /////////
      input              TD_CLK27,
      input      [7:0]  TD_DATA,
      input             TD_HS,
      output             TD_RESET_N,
      input             TD_VS,

      ///////// VGA /////////
      output      [7:0]  VGA_B,
      output             VGA_BLANK_N,
      output             VGA_CLK,
      output      [7:0]  VGA_G,
      output             VGA_HS,
      output      [7:0]  VGA_R,
      output             VGA_SYNC_N,
      output             VGA_VS
);



//=======================================================
//  Structural coding
//=======================================================

audio_nios u0(

		.clk_clk                                (CLOCK_50),                            //                         clk.clk
		.pll_sdam_clk                           (DRAM_CLK),                       //                    pll_sdam.clk
		
		.leds_export   (LEDR),   //  leds.export
		.reset_reset_n (KEY[0]),   
		.hex210_export ({HEX2, HEX1, HEX0}), // hex210.export
		//.hex543_export ({HEX5, HEX4, HEX3}),  // hex543.export
		.wifi_RXD      	(GPIO_1[29]),      						//  wifi.RXD
		.wifi_TXD      	(GPIO_1[35]),       						//  wifi.TXD
		
		.key_export    (KEY),     //    key.export
		
		.i2c_scl_external_connection_export     (FPGA_I2C_SCLK), // i2c_scl_external_connection.export
		.i2c_sda_external_connection_export     (FPGA_I2C_SDAT), // i2c_sda_external_connection.export
		
		.audio_conduit_end_XCK                  (AUD_XCK),              //           audio_conduit_end.XCK
		.audio_conduit_end_ADCDAT               (AUD_ADCDAT),           //                            .ADCDAT
		.audio_conduit_end_ADCLRC               (AUD_ADCLRCK),           //                            .ADCLRC
		.audio_conduit_end_DACDAT               (AUD_DACDAT),           //                            .DACDAT
		.audio_conduit_end_DACLRC               (AUD_DACLRCK),           //                            .DACLRC
		.audio_conduit_end_BCLK                 (AUD_BCLK),             //                            .BCLK

		.sdram_wire_addr                        (DRAM_ADDR),                    //                  sdram_wire.addr
		.sdram_wire_ba                          (DRAM_BA),                      //                            .ba
		.sdram_wire_cas_n                       (DRAM_CAS_N),                   //                            .cas_n
		.sdram_wire_cke                         (DRAM_CKE),                     //                            .cke
		.sdram_wire_cs_n                        (DRAM_CS_N),                    //                            .cs_n
		.sdram_wire_dq                          (DRAM_DQ),                      //                            .dq
		.sdram_wire_dqm                         ({DRAM_UDQM,DRAM_LDQM}),                     //                            .dqm
		.sdram_wire_ras_n                       (DRAM_RAS_N),                   //                            .ras_n
		.sdram_wire_we_n                        (DRAM_WE_N)                    //                            .we_n
		
	);
	

endmodule
